package param_pkg;

    parameter DATA_WIDTH = 24;
	parameter MAX_DATA = (1 << DATA_WIDTH) - 1;

endpackage